library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- Entidade principal do sistema de m�dia aritm�tica
entity media_aritmetica is
    Port (
        clk            : in  STD_LOGIC;         -- Sinal de clock do sistema
        reset          : in  STD_LOGIC;         -- Sinal de reset (ativo alto)
		  ok             : in  STD_LOGIC;         -- Sinal para fazer o calculo
        entrada_Y      : in  STD_LOGIC_VECTOR(15 downto 0);  -- Valor Y de entrada via chaves
        led_resultado  : out STD_LOGIC  ;         -- LED que indica resultado pronto
		  s_reset        : out STD_LOGIC  ;         -- LED reset
		  saida_Y        : out  STD_LOGIC_VECTOR(15 downto 0) 
    );
end media_aritmetica;

architecture comportamental of media_aritmetica is
    -- Constante X: valor fixo para o c�lculo )
    constant VALOR_X : std_logic_vector(15 downto 0) := "0010011011010111"; --9943
    
    -- Defini��o dos estados da m�quina de estados finitas (FSM)
    type tipo_estado is (
        REINICIAR,        -- Estado inicial/reset
        LER_ENTRADA,      -- Estado de leitura do valor Y
        CALCULAR_MEDIA,   -- Estado de c�lculo da m�dia
        EXIBIR_RESULTADO  -- Estado final (resultado pronto)
    );
    
    signal estado : tipo_estado := REINICIAR;  -- Registrador de estado atual
    
    -- Sinais para armazenamento de valores
    signal registro_Y : std_logic_vector(15 downto 0) := (others => '0');      -- Registra o valor Y
    signal registro_media : std_logic_vector(15 downto 0) := (others => '0');  -- Armazena o resultado
    
begin
 

    -- Processo principal: M�quina de estados finitas (FSM)
    process(clk, reset)
    begin
        if reset = '1' then
            -- Reset do sistema
            estado <= REINICIAR;
            registro_Y <= (others => '0');
            registro_media <= (others => '0');
            led_resultado <= '0';  -- LED apagado
				saida_Y <= VALOR_X;
				s_reset <= reset;
            
        elsif (clk'event and clk = '1') then
		  s_reset <= '0';
		  led_resultado <= '0';  -- LED apagado
            -- L�gica de transi��o de estados
            case estado is
                when REINICIAR =>
                    -- Estado inicial ap�s reset
						  saida_Y <= VALOR_X;
						  registro_media <= (others => '0');
                    estado <= LER_ENTRADA;  -- Transi��o para pr�ximo estado
                    
                when LER_ENTRADA =>
                     if (ok ='1') then
                        registro_Y <= entrada_Y;
								saida_Y <= entrada_Y;
                        estado <= CALCULAR_MEDIA;  -- Avan�a para c�lculo
							else
							estado <= LER_ENTRADA;  -- fica no mesmo estado
							saida_Y <= (others => '0');
                    end if;
						  
                when CALCULAR_MEDIA =>
                    -- Estado de c�lculo da m�dia
                    -- M�dia = (X + Y)/2 (implementado com deslocamento)
                    registro_media <= std_logic_vector(
                        shift_right(unsigned(VALOR_X) + unsigned(registro_Y), 1));
                    estado <= EXIBIR_RESULTADO;  -- Avan�a para estado final
                    
                when EXIBIR_RESULTADO =>
                    -- Estado final: resultado pronto
                    led_resultado <= '1';  -- Acende LED indicador
                    saida_Y <= registro_media;  
						  estado <= REINICIAR; 
            end case;
        end if;
    end process;
end comportamental;